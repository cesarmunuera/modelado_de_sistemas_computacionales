
library ieee;
use ieee.std_logic_1164.all;

entity teclado is
  generic (
    REBTIME   :     time;               -- Tiempo de duraci�n de un rebote.
    M         :     integer );          -- N� de rebotes
  port( TECLA : in  std_logic_vector(3 downto 0);
        COL   : in  std_logic_vector(3 downto 0);
        ROW   : out std_logic_vector(3 downto 0));
end teclado;
--codigo inicio encriptaci�n
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling="delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
TnNtGfvGGbpz834i4y37fsq7Jv0q9cXV19mJsn8VzYhFtdwBsVzUXbrgY2XJMXhyxOVtdLA8jQyw
T/ZLJwlOAvsVWmo5qt1xVQYE6JKEwbdgVMKOL89wcdRPDrks9GERsW2q1hq/duF6X4Gak0kg+XQz
aMX6nS7QImAYQRSbnN0ag2lAMQGtXq6l4HwFJcG0NsPyTWTBQm9OQxkCOWHHX50lPRmr5ZVqB3rV
LOVK3ObzuXNWqGohHei+QeCQ+FnpWYr5l2qQ9mKI7myrOdM4xqPH0l1cXxmuei3vUtHthj6Gqb0Z
HK7HrJVbqIx4brS5+NR9MmDLbWdfRpz+a+qsyQ==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="IgYwHDyVaG6jodDCM30HmtbYNcufjjdhuBpHPBPT4uI="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4208)
`protect data_block
6DEZY6WzxDSCk6PE9HWRWvXrfkgPKDUx/ndrcGrOfwNpjs6K+bLQEurlrCA2X85xAbWpFcaQ3W24
doeEA3nWdGxr37wDqCkrx1mpfovRXkQf6CHK40GoQZ4iEN0XMSynsPSY0/LohzBaWoBpeSSi6R9u
Gcaov45xoeNaF77Tu5tZjaY335xXyuDP8dsfKoEy3DYaIjsBo2iMiStGeTes5z8BIXKx1VdyN2tz
Q0VU/G+ojmHItE5h+OSzyg1js3AUzXoxoSZWkfgc8tpxDdP3PLKM45XQHJA5lpFw8lxukNYEAqSU
3KU6sJEX7uF4d3DQxQ7URgL3LRXIQsujzd4VEWneqSpd6Gnld74GnXS04OIRFIZz+i+z+tJ3TADc
teeKkFTz1+OAAmq5PbUfetLlN2DgbYVHMDujXisSkxph+Ac9ho6Y9k9EUt6L5GIlBVUpt/84IYwK
0gh04WLAVoEuDUWPdMdLFkt4T1iO3VDPfpvDx/ghmnwV/2y2GyK+hyh8OAPQclRRRNVHhPEhfEBU
7/tvAW3yiXpxcU4gvvEDPiS5eJxQBnNCeiRMDV4CvAfcXg1dE4z50ZxLIO8dq+X0lnmQTyTwEv++
icxN1lEvbXIhR4ZPuU5iNRqtM82o8ClIk3dxISkOU7jfEEAITRG8c34qVMNHI/1KjrmiqZAFpBPE
uqda8uPNZZIbI0YMADBQUXnsG5822TOMOE47UdBs4Eutyp2RyZKLRD6i8nxdP2aCiqSFDiIxp2zp
XzO/AKU3nCV0tO4ie8qPS76yy+0+fcpM36PE9MCgtvnoyJbOGB5YUpVxbJnUh40ggDPulrxl4JFk
XyyQBXzVsPc7m0Ls0e9TU6Uze7fwEXHpvk95RW58plaVSpZtS0rpe4kSolsXQs2XxP7/6RjHFgPE
w4yhulmZWKDzM3eNVRVubEhL3V2uEEkXSXwgMsheS/d5ImLlTwG8/jPxgD6jootbQvdp6vjqTg3u
yUc6OblrqnRC73frhErYLsvlfyNDz2x3chPlvFBXaXf7ytDCS8JFfwqs6gLSW+EnxwXAaKZnlOB4
/UEV06Uzj0x6yvIo/9CgCGThDAXjwdFOfimDWwSXWbIy/FsJUYGB+Y6poaRhVLXHdfIkUyACQ2Jk
YvOaccyngMvYslHFntQxYR7j7q+uBbcU1CpO0ezbVgGBUkOahLcd3/TS8QeiV/BBimHF9nMiKEKB
rO4V4APbXmHXXcFieMth3FbndB2lmbQ5VcJdJXlttEGQSvs3C7v7YjeC8jYF9S+PMSDKWpooNtoe
RUGtBlMGxyLRb6QPEp+k7aZw3qqss9+gRm6kMqAOG90mCWnpnwh6B6A+BIk3VICSy+oE/Dja6VSr
7STDIsxZnhIMQtVop/1r3M+qBEoXPLnwkpGtUjOvIFQTYqz7lHpT95vLB7h19zWUH6x9GhClSzc8
fgc6PHfi0Im53NpXXlynVokMiP1cJMj66uTKgx47uUt9r4QkduSIiTAid6O1deyFIBz76HS9xZbF
afyQr690PdiD/nq3yStSGv4K4d0T5VK+KxVcDzIq82etIpGVSL5lAlYHXIujO5HtXqhqpJoPEnbK
WMQIGS1S99gqKGjx3g2A950/hcPcJffXnt5bN7/JBqkH043fnO5nqH6OGWY21piLnB4hGuAd3POb
e4ooQA9+VADdCZSa5IctqYHuvgfG20EFx5Ui8nGogle18w59wA55x9ruVhhLefjucsMKKw6bzAbK
yXU5mpnhA4MHXMkQmJXurdg6dtjI69mjK7P7FCQljvu2Jr8oKVlinJfWj+jl2TQlGl+FIYyF1+Yc
gK+ya+A95Y2cpCyD2tEhIgUmUERbKqBHiyLVGl9iUkmhWAvngxwe1k94Z5kG6q6BmNgfdVfAXeeB
LuxeDswPRBiNtTjpOH4I7XMgWKIYB5MEMZ7fWXnPDW95fsw/PIweAfXF3Am3GeB+WGHOesub7Kf2
R0xd6Zv+KEtccE2S+FHkPBn6ovIy3sXdL0xItWR9yOq/ivbp+YTzXrmwN/HmWpnaoJS95gES/eDH
X/BemuCcNiM46lU6Jf7DNZZPbXnNQnxqedexI1IlJuzaTQW1KQQXxKb+JKg/lR1Bx29k3l6dk58e
TU7m+xi1Ngf+5+Ev9FRwO0tpEM6sA4hX2c+7KmNa8Q+yQQlpcDkXYIzUGBrKEgZYf+2vBUwCpNA+
H/2sq5oirqd9v5QkZpksDVurtW5pp6PC38Rg0FxIX2E0dCFO156MyCJFZAUayYiS6AomHr7w378t
RFzgMmfuQn7/YH4VRcJTm83LPPWuXqZB/sTsY6BWeGVQeNLUh+bb3hVIjWr74jTaWHnyjttA/syZ
Lx8fS9+Fh9svxOPpOWjOs1nRxZfX8agnlu5BfcAqYwzeAjHDEhIaAQwH+wUfXrLa8o1EUyvbGhdW
qGTmaimPcaM71P3s2DHwVjzIlI8sL3OsdqDvfNoDgGVM5T/Aq124YP/LT6tH1fqy5xUohaYdVtxy
THnzNLCNH9BaOyrtWD63d+5inZONB/jjwjmbu1IC9xHfND2sq+knWQHvKQWPAw/JPGS2rwvQzDWZ
/1C8pYRy9aEulzCpgQ2yepSin2Piskf2UOLFmFnGjsxKR9Z12893Kf3Hba9+Aw4w5s8Njb23T8Zw
nyjBnB+KZxcNoFJNmcbgu0mIA+RewusJ2Q/xWFgc2NAi5vnW0yXruAgee3YPFX9yNQTxko88lUOC
FDPuQjrSiynmXhabAYttTIF8f28mblWgS9WOwmqcYi5Mbs0QAOTEeR0sGU8ykYZzaY+GCCozWZI/
BU/6aFCMg7zXUcKnB4JhTeukpj9QlwJJ0j2j7hI5Oq1pt0FkZvTqfZN0SLG4M41tNTZZhdsaDs0d
GI3cdNNeUwSmdLbqbCnRRhJ6jWVv8NqlEaqMFEV3hWFEcoXmOFmhwACOv64XRKm9a0S8e0R4aKyB
Z/0Yre0Gtmt3fk0pj9iHRyOfQ/Kd3g2PFme9/gxkoILRl374XJ+GvUts9fUMWQQ8sgoKWteYDLNC
ko/4bh4hFCouPxoCaetchOhR0taT1M9qqeAmeVaYs2dsjtz51AjGrOVzymn2p1pmiQQpQWn1YJ4L
UnWDnshNDi0z6Qe/ZuDcYUMFPClqGD43MRae5KghqEQUdgHq2qO8Ooysl+sl7XW4kk8fxCVVC8Gr
KlG9Y3J8iRRxdJcTOrPs9PadKdJa6HuoBp5MAtRKa5WW0DQ7IgT3rSK6hWBBB4QuEizc2/Z+Hv7G
V8/6S4MLF53bEzKd5VmkgWGl3I9kCGU5A5H1LofsfKTA/IYbZPtZbDhusPklBXFEPte5ZW/eDFsJ
SVYwjA5d7y65KVS9n8o5eCIPNbIidmaLsxCmBC71o/dex/DcBwk1GWJLDERW52pv80KwhCTlp7bM
gKhZYU6yCEvZbGDQoW4xRRgLDFsYU7Ois4HOWAUB8X16bPgGr4mv1afkDDiYBv5geTMcJd+u2FQG
lYa0JaLTura3w4wY4mkMYyj+nFLiDgyu/n34FLRDqNYpWxCR+LQ2M2XvbJMIKJOR6iMKW7izDHy5
jtaWb4p8eb/9tmKMArbMp7iLzmw5WOMPjhUrYCj5uJOoXrH235hjrX/cIm+TuAkmANpYI28gAyEX
X4x15mwj52UKONbQzfIAaTP+6JBB0WKs/qPeQhJEJrkhSTxTjr05ZMfajiPy2o0KX9VxHNkqXLBN
VTxLRZXYZM9Y4kjSh/OEMVIJNcx7vgX7NecpchjBm753dr0ovaMTSz5z1NnXMX8jaGI4u7ZvrU4C
rKpmOGZLuBaR96LohzAQkgIL1zZUQUjLGoKMPiLUfvp+FJeEH6+d93YvJUiS+ZJxjRJg5/ulZuKJ
ZsPPq6dYHbfYgorKxXjph4qdM2R83s6JBrDf06egS+imHok0zMlzRBLgeCgxYWFsoDXIP609zGn+
BI8BTnwIbTpFH1Hx6MR4QCe0GgxEYW/QYOSWWoUD3aUiC1F5UDLtoS2pm77KgPYDnXs02sa+GE6m
20b3Zg43MM4ku7Suz9tZo4ybaHxE0w+GDQAzu7jdo34yjZQC3QUeG3XbsLGE6QIq3TWMU8zYL1Q+
5Sf8Ic3Fv12UQK6sdKaU/zq/rpElmVkFd8ExypMr+TsZYhKZCG/7DDe9WWIWoXLq+HVlIcUiIz0M
2yy+gmpvwYACRDNbhNE0TPANI75q6TcluID1uRkqR6D/Mu8g77WK7qgSIN7jxu/XgOMQ0E8xur2u
0Q2PM5d5o1eZkbn98G2pYkSeDRnuF1T3TJjgxAk37zm0r4Tm4VyfgScqRZQ8hsYX7z8HiQJvMjgg
D6uXZoGxfFi0Ga9/u/Jk5I/M10Ol1LpymRZhpBFzRx3qzFPf2w9QKuEID54sCcmjQRGPBUc5+EV6
qJpOUgAZHAW79Ws4UEYWb+YC7FFYil6kgHDtxbKS1C8qSubpUskZY5wQSeAf7lQoETsPgyJix5cx
ToeWN7+BbIJEOb+6lfCd7w4lro48q7YW62oN4mnDLhOLQ7NdQFbK6I9HW/XqJphys3bzxvKWRSNY
PbWVVSuVahiFw5ASV+VatEJ+gNMGs3DgoKfeL97lBeTnAujYAAzoiR1QIDp+H2WS7cYuk3kHOAaa
T5iOtWt8yHoIbSGK/+cqdYzbWIpQ4GkdiLXXCqSdRs+C0NQ94dVqOqyz4YYpnrPr7Ft6UhQgFS7A
sVcEzyGNLThI4PyI+LQnUE58ppO6OCYsDzMe+oQBDdFIpfapCRqxpzheQxy0HDIANlh1m5/adsl5
BlPX4NdAQ534NCF/XwtA/CUI2kJDceGkDTA4gwvp3hq5M/I3TQtXqF3V6iKfq8Frz/O51gQirqlE
gaCpHoeETBgreo1b1Ilt66EaUGs2S80LMENBh2l3iU/0LRyBBvXzIIDV1uuKgl3WhRPWInRF7+GN
WBal/hjWAz+WDRI7AXi9OZh80vrlh3dbusrId8Hok9o2OuvSURZgL9QoWz1pIoyglwmYcwWgi4Te
tLmgwrR17VqbgZlZteh1h03BbS5yZnUn/RyJI/HhqyglrrV27Cv9eEBxTNYmMYb8v/9VLy3BhTRJ
LsAKRpQuC/msNO8vKAxbB2lYCHkO77xAESbrqVD1+TsSqfSu4kvF32ULl5RNEgDbYoEroFMyyxik
CWmghPqHKR3qmEqHiSLs3UhLtJJh/J6Tbs/lurDK7pjlzB6454XoV9lcDVhVr6KImHcNARzxC9Pw
127ou6vnVz723Ereqim0q6b94+oxiIxqdavcYXew85w8NjuxNyYmxzuDtlspRe2dWl+QO22wUdT6
gcg4MflcbLZtPmdGfyUV8QWq6VUSUFzjUslN5Aw3vqNCvbhlqC4QxOcXT+VwdEPa6tcFes+KIfOT
B9E4DhhSqpMZMPMuZaqXiHjCsoVWe40ipCVb3jLNn1FJkHip8+s/i8gp/39cnApE9ehy2yIRIKka
HedGP+OVXtRLfzefZJvmMgGHZQgw0vOhmY9uJXMjj7s977U6r3wB3184no5yYUrueW83hXTzI/bO
zNp5IZ5KvhXnGhIhE0lqcJ14XBST5cn8Oeq3GqVO/hUWx1/Rk7+QcNIp9vFnysw=
`protect end_protected
