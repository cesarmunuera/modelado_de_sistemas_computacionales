library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


entity oled_controller is
  port ( CLK         : in  std_logic;
         RST         : in  std_logic;
         DATA_OK     : in  std_logic;
         DATA        : in  std_logic_vector (7 downto 0);
         DATA_SPI_OK : out std_logic;
         DATA_SPI    : out std_logic_vector (8 downto 0);
         END_SPI     : in  std_logic;
         BUSY        : out std_logic;
         RES         : out std_logic;
         VBAT        : out std_logic;
         VDD         : out std_logic);
end oled_controller;
--codigo inicio  encriptaci�n
`protect begin_protected
`protect version = 2
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect begin_commonblock
`protect control error_handling="delegated"
`protect end_commonblock
`protect begin_toolblock
`protect rights_digest_method="sha256"
`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2017_05", key_method = "rsa", key_block
UgJM2jfUgphriBqjp32zS6HYkSbO0qbuRJaYfJhJgEHPGTgtnyIo6BzIt4PuGS88+4kzK798M4d9
OENEYYhXRVsw63M4yYkmQkQyhKfgEFrnAIOrrI+n3OjFadQEmAhbZDJN0EzBJm1NfiE9hvSNUdSh
xSLCYhhFp2NOcasCQZvBJiJD2eYZNYd2z+p88dvBy+E8q6F+Ua+GpcbwuL9YR2F0/KbdTXbyWRc4
Ps6G+OHLl/csS1rKi0Nh+d9t3TC9sY4C7sgxgBO1ybUEMkevCjfcaKPFC/bzLtju9/wk2bUFxgkX
6XBZyFvaKEXwQpPTGIgJGvvX1WdN+CMxGEmYEw==

`protect control xilinx_configuration_visible = "false"
`protect control xilinx_enable_modification = "false"
`protect control xilinx_enable_probing = "false"
`protect end_toolblock="7FEhTe2BeZNo4AbR5JLL5yzcT9c2phtgKocAghpNRhA="
`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 21568)
`protect data_block
KiWTsmVNXw2AGjrN/2qDJNMtPe1Gr4d+zDcoX6TamHMPahiqs4MpQZ46SIBu2A5JyHv1nNEjUmHt
DOISJTmOwvX0UMtYvfT1SOKbObw3co1I+EjdPW58zpSdB9LwCVcYRmX51w5LCuH+hr9DonVNvaI2
zrURoe+E5BMl1R63Q/I4FqUO7/kOO6ZphqrHe+E7KE1IGtzykIzFmDntoTUrVkWz4oVNK+fLgtAm
93Zj5+YUKOZN8vG4ID4jmSa8DpqPs019LcnefhKJ8K8EmOFvz3MuQFesZaWR1o4V1izz/BrkIAxt
wNctG/xHtiVlqzDAek+v793t5GP1tyTrIoT0pjODesfcZ370umEnqmDAm0gR5ugv8F6u64jHuqx4
XcPnU/p+TDTJJ12HbAKzEwNxscsE0x3h2RLVGmVcXUdKFhnj6n4tAhr1SMHM3pDHMhBYtMV8GF2u
GqNtpLgF6lDXcNVp+fxtEl0R8KqcrVOpqT0gIkIY1r+0MFB7xytvUsljsM4i4oWEsrElGxd+LM1w
7s/3ch0gIxdaW32b5V6aiMxItj4GWNN89UjFoEiPBtf3tEV0Tk5Y4NpIx+jkKdezhGYJNUQ5h6J7
RHOI7mK/qcvfF0cO8XmsGqhaEMDWeVBxJ7lyiaqj0erMZ5OOwitcMlVYkWqG55HYAEkgSFKx8IIY
kW8mHvUzGfH5yIOxwzHBpiQwL87+aAGCVqY97QHB1m7QpDXOTwtEgXUCHrK2d3aWikG6q9LWJpQf
JZSLR6oXNShRpbL1o0nCU2WVRzZ6Z1ln8L+tMXMfHIQ3fWqlSclj7SAHrCla7T60dGeMlegvFLq9
TVI2Jj+Q6ExrBSh93gr6MYCRkBs8RxphQnhxoAKNu3q3B2Co9S6e4bm/gyfCJVzT9EnlBBwfG4zw
qSFWK23LEl9cDtKjXXelaMG6WaCWmqiuddu7rfPuXbDuHWxnWC++7UnFhScK5eK0wXr/qorfbDup
qA/ILuGa6wJ2dpv0yL43Yv5+AQ+16zMsM4YNek3VKMsVI/fP8/vkN3wKOSv0FOvlRoCWf8LAeVaQ
u06In2RFxX+h21Uzk2KvEHPz+2NaNCCqWhLnAuzCSGuZrgCj8b4LUWZf006do/n4Is6Af+WQtykj
c/eU/dEqtNjiWtCpCME7FqzXK6FFtAEdr8nk/BB8glOKnpT4bDU8rJT33vgRKwVSSJ5tmPbJJb0b
gbyHOlfOxU5+Vcv4WP1Bf+hoaN2w0WpgG83yxliEQjeNN99NU3MGZKrATfac4UJE9+xJbTW915nc
PJqVNWR1i/yKL0GWEnQoiOf+aD+TPrCiX7AJZilyfm2yO38phdPX2+t072GBEQDkPpPDgQ1qDfbg
w7xUkDKLN7urnbcZ1RaztAWehqfhcky3sjt5Ux8oe0lb7+ch93ik6k5QZjTlt5cRpDO/I2ByUXZk
OcU/EJobjVxrhfUByZFje7HULAJgwgeFovC+Qwys/vNE3kiiKbjWckeZtkYtEmtq+P1R5Y0Rq5KO
8Gh6YB4SW9wR+4B6cSmdJLphixqw6bmpVWNZh5RV/ZlfzqVpKKlQWX7wYn37KNW+HcDBm9FWSSGJ
ijQv4WFFYTpomEGURUJthkVLmAe3wVBJyQ81RrYCI+GQKtaLDk8wtywKQ3/cXUehmGAu9/kFumZf
83p/2be5Plq844MvZle3bvqV6L8xOD5qZmoa7V9z61YqmwRou/p6LlXZ+XYSD7NswxBwa8WmcSDk
Acrlo8Aw5L9meZ6X8xoCnum1w/y+oftw5stK0mFRHlryAvNdfbdcq9a/bE3pUS8k8ypqEl5Yaigo
S2cEUDBj1c8xQwa+Kw5UEWJZWeA91Geb3aTWcFaOamGohp/6UnWCOgSJKz09xQdCGJUBpEsfRWKW
s6uK7oZFFRyfuu9Ad6ZxQI6AReb1lSzYLloRxLWuL4UH+2fC2Dp6k/jGxSw17C1QGgmLk0syh7JZ
F+SLTjuduZjfj+ZeN6QhT+zObD3KUiVw3xcy+pe09ukZG+bpAxTymTAykv5jgF7TnyDEZQaqeYbv
AI7f7jcb3ihaUOjdw8j7UA4sOFGIasLt47XzROiU8Sh3IwNae5rZunhRFwz+NLIws03+xpSTkL47
AS1NLpRlUpqw2ArKWQ7MWu2T4HA40HLzNiiXJzos/E5REqCuF4i/eEC6R17fLhVKrkdd98GGQmF5
+v+kWctUb23s57bYVdP+ZxZyE5ql8NfQS3cbRkBrBEh4nDFA8RKazaHJsoFLbI5g/P6JtOMhSAi8
O8VkkPTlSjal/9VdMm5vGNqwhdF+0qNUnAufq9izut3EaQd0W6dK482TE/pII3IzbVXdPuNGKMaA
Q2fenl17N/EG70z2QInyfFc8svbrEDayhmXljYf+bJKGGkHgKM5+NvsE3KxNhTPEaRT3GACO1Tmu
dMFKsVRcR8bpy2LwOIR6rZ5KP8H0QJtTdUO1Z3gDT06kZ0g+nZ6S3/8uHVer1KWfgsgyHyaTzCVi
QZ+XI9iKm2aP7gG1otBEbg+mOxO3QxcowNjJ9tcP4qM1HPoaCpr1FP/FqSx66zAE5wKhMa3z+SBD
8WNR15Ji+A76BpQelaJZu49r5VH9zlMeRNYdzUl9lXM+dpuV/4bEcTpTaH6PUJgqu+UC+KHbJ7Nx
SLqmMTV09eCEssF2xMSgOsla+abr9cPtZ5fb/cevMQMQ+vTzP8runDZH8f9pmFkyvPCzXw3YmH4U
2ZGxwgI2T6J/1/kGZmNru1AmnFiR2PjXueFCzuY56M4Hvx/GWyfV+cR2+hlbOeBvSgtFxQZ/l7op
1tBUyJqqx7cEt0Ogfnaa5+RImFdHXXAT1MMwfqRDY/Sz1PdHIx6D7AqtxLSdwRoh8G5I+WHOkEiq
dI49L0Pk1no17aEwoalqoJ1BRVCF69dlBWyTEoM5XYv4UrBzgfRWBv4x+IF5SwDHoEFIDWL4AgTr
YzvHxqg6J4v6ZfRSLOmoYtWT6eh9LvVY6Diz4c0+fIOiNKJ2tTz4zXc8JSFgEuk76KBcMvTKexVh
TcfHQn9nnIF12uFv1PX2C/wJLUWcpiKUKn6BDDj75IdljXNbxguM6aF0SDjlqL8dKbYtV76rJDyB
PrtFpN0q34QmdBieT35u0OUphpQmBO2/JqrM/nTSGndXuNuaEGsh5Z8Js/SKh2FULdNhLSsAJDq5
12Us2Unx5zafWJclr6lblNQK2PRoqiHe4oZrDZIUUfUrYOcNgEk4iXAEQHbMgRHJgDgblLgcdpGF
bJVc9ruHKI6jeEpDHAnBJUlcc0N8ns62JSfRUEMEMzigZzaqntspamm3Y62hNlzLlv2k/SZmorY2
LUnXl+WDXDyv44dSLZGoeaSffZJNWSkqzJqP3V+jbRLZWoC5V+n6bYbIL+R/Tm69suNYzH7ryLXc
oB5ga1jHHGbQ6v4V7VzFaHaio77lBGfau4fbcdejbxojDFv4MPGgIjIgjzqcWruc+9zBlya/fijr
HgZbPwq6n0rg7UNnRWX4lLFXGqGCyW+8JzN0MC4I+V34RNm9Z0hOPPznDkEm2CvxUrtXZTrM2tIH
wZQDKFjKxdHmeXt07fdKXcbp4yN6jRQzFRKVpnlKIM+vGTjHZNIzthIm+fjnArZZeJWdDYlbmFWP
jJHeays3O8F/6q5APRJsXKhx8tqzV3BWpk2C9IQt+hzwboucF5eIRnqekscZry2kn1QBs5OdoqMD
JU48NIPAcnd7+fKLs0vuvTzWt1G5bTXVtsiOXfbOd3JQbZzGB5xBQ1b7bZ3oX3dbwXwSD5biQvq7
nggfPgyZvRyo3jmrVfhnadhFStMfzI1uFDKbS4wMyW3cJ254S2aCM1QRapVupx5H37A/xfdq7zYf
nQFNBE/TcAM8uxwQ68q9cEDaG9yGo2o4WBOSk2zDLNFkoi3ZNc1G5SgguegKMax5uEL8wS5ldpX5
A/r+5fWkoW8gU6F6P2pSEmYjWu0dDt9PKHX0hGHHIruKvBLoY+1YiE+OiK0iK/DlJA5K6ca3kLnA
UaeYgh87RLogUgcVy64cCoFgwlpitb4AkwcPw1uvBGs6xVYSCeoYD4/4jmpFmpyZfmSNsYo8KJn+
sbdhH2lSPs+W6tBa81tDw0lbkEoIbsFJN8GKRLTldsBWOcrODxxIab3lgaQ8XUEFB6aonf5H+OoT
PwYpX/JRfSlt6I5okZuWogIotmM0H/EJa9Nv9DRU+GFu+ZvGq8Efx6wiMu99FCHe5getIfluasa0
AgOlwOoZ5DT/Z+JEEcBK9fTWlhocfnXIgG03RJfpz3gtOzwP44MAeih8FNoZkfDORTGT6JuHCEXD
noAcJ5kujCi23Z4gblux1EoX5MtxiEQxbLD1WZypS/l0z9zOwSEi3Ufg58cvW3wL84ZmHE/rFdVN
yTLJCW0bblxZg/tlW9SKHYZnN3ndSUHc4M5ZTtjopgqh03mq9+jjUj6YRnz8UtX7nzufzgdT8Be3
xJ1W7BmUB4t1kk83N+0l3Pq3qvYWnaC6g/swwGLyg90gnfT/gLHc3GCoWkw5yp/Epka4lHUFmGOE
S3bQ8LmkKzKFKOv2d23VYcxBCjG05aGu/lPU5ZFiP7VTJcabWaqYmWJZWCsTXy/PHceXmER8YGHP
HJYNvMrUoUhxOAid+6kvuI+kqCOP2NMFJ5//LIsobAlNcD16Ugzbhc24Y+puwJBzNWVDgjt3Km6c
i3g7XWtst8F1ZyjJFy9eE5Qu35Q6X65ri44YFnj9CyHu/+0DZh2vvG57V/648O9308YgZrd0fbir
SAiFCC+cH4qhSPyIKNTcGtMawe49XWbccxkTd9JiURSDx7MeoCGdUtWHK0SMTbaBDfI0WPqk+X0B
rId8fUkrPMdA3rQH3TD03Ciwmd6m0eFUD5aZdeFdjoNqvdeVv/4TWviMENMAFem+t1dQGbJ/UWhA
HxxLiww9vDXodBFugIBBBWdNbSRJRguHNp3GlrSQmzQBQv60GZvkfEbIuwwOwy1AUv0ze+uuqVZ0
wOHrV9nGVgiGjoR6y4Jj55wx72HZdenTs5FBH1ngAGO/3ZHBBPyCUVtK5zAxKolcrgUrGY2yp2gR
8qOIXrj8uEpkyeYTw98DY+ZZ6xiF2uzBGRph/Qldi3qA08IHZdVjP0PCfECwgnV5MXgWDtpGvGAb
6CesQV3/FJgHR96mIV1c90cZTQGwFUTruc9m/dUtTvbaXIYzVlK+PR70z+oODoTrbmyaY0x966+e
v1PW25az5l47T4DZmw63obKUoFcWjS9cITsU0Na8OriazJ6u+u0a2lsVo+PxTfAuNHU4Llx1M778
JhXqTWsVo2TybUGimSw8PFobP4b6X1fSFsq1bll4T46cz0Sb8RV+Y80/Ppt1OMLRiVHhskZWsFh4
/F16UWcJx5PAytx1ClD2aTpVAgSKOUcYf1XCAc7WfWv5yEyTFmPLurLlGvUWdqV4B1NgreT38YWY
YY7oSuSsFqNJJJWXaynxXSkgukGJ4sOBw+/0oCFNY+nCOEazg/ghFnCDGvSUw/RQMgTuLwjUtQqu
yNYIeHj6ciuOlWxT5j29Ypm/S3dYhREqf5rKOqEYnEcuzIPGQ7alCoEP5SReD47wZsLcLyD+R6RR
m5GaUoIP9L7POlI+uBfkNRcMvWb4m+a874Xgt5+datGxNw3D69WDc27Bqow7VfqlCtjpMYMiOsT3
wXObOs5uYWHJKe3X+loIs/DSxUZfWEFPCtupaGEAQwfbobFhR07MoB5D3QX1S+x83LyX/6Cy78oF
LzU5766dZnKejIICvKRjlC/Q8YV1C+ozWeh/qY65XGXybHTN3zexWd2xXKhsSG4eS9lGT+hmRBJ8
X8rfK0Rzpk3oMHDzAVbT1NDU5nfb9HoFCWyb4RdCvkSZoybQ9ANSq9B5+dU37sS/uRmq3QnH4hXN
qsOWV/wQFH6o89GU2kiq3XJA8oBF2MUmloh5Rb6MopmQqlkK8atPGPalIrFLSZba+bkKknZjGbCt
qk14M7cNFGF/HSRoz/2DkhPRvvoptq+9sZv4M+6Ci7ViD6xSuD6H+7DOPgcvDbXBpXT6yPDKR2Og
CWnXdJZ+78PAxkDToG/fjmjYHjxJplgS4BAGCBMOldT0XR9LvlNQWEGfp4quwyXqdjn66XXn2QCA
nFolUBvQkcub+nvPX7uJoPeirhCKcX5q/GJgSP3XvgtSrty56VaOl9BXGDwvK7v1o91kL+946fjb
sgoePBNHi2xVIll3GL2z182QAhtS1mEfYd5euc7kYBrfdo8T9Xkx721CPf8/8RSLFr/gxiBWTvmv
rtyujFYwSAC1AnCAJcqWGqYtlT8/kpRS8yxpTo/pGD7tt9MYBvD0MW++/ApJ8LzAh7nnit+RJk0k
kf9P+gqEGvnnaxNLf14qFlp3qc1uB5mwRtFnB/Ny/zVMW6qa4geUD3+cGhoo8WT7Vu7pb7k3Kb7w
GobSLYZGo/L4SviCg+NhaXoN1Iu7EDnWGtbBeKmwgXXmI/rjnIr8bOSjriHjZ5W/eWwPAbJkUJOq
nxlKae1oufFqt6q+Cbh32/RfXojQ9Su1ewCYG8R++kMUK5tk3HD/TQX72jviZwaMxzBspYDD8MXr
Ab82hwC8QYdSTNwq5tPAqGoaCDhnxV/ocl6BjFhYfR65FcijHx2dJhAXSjn1a6jVuQus+FQNo8Co
95AbmrAAvmCO6nZ6uIOBv2xVA3x9QmrGTwGoR17AQ7V4xHKHBb3QZ81DNSt/+IU+lpt53jcUGqyv
766wOydQisIM8sqVce++1T8HmuU8MgKXKkTSawe0LJaqr4tiEbFBtGA8S2PPw4FRyBFt4NlPDkrY
0B3gcGS16gKho39iL96dkyYHgYAS82zunY5cDVyND07pcniPkucgkT7juOjJGk3AkPfj3A1CLYAd
xseOhZpFOumLGpzh0FHPpSw91NT8Jjy4xCUM8upw73v6iCEdrJyhlocGWQVvP+uAlptUfoWIUTPT
3Xu7/YpHYglXQvgtOCOdOwd0XVhVCy3UIt9U/dZ7YX+wNR7yYCvnZvbEepEXZTfNTEQesScxwkEd
+VaAqTJowSuc3IHzI7gA/MDWCn+Y88QkKqnikq7UAGgc4A36NaKpevrlztp5pnLgynl771zLHG+6
Yt4TsxesH56dDzVWp2f+dXy+RjncfRs62hGFXhV9i3kGagXU0U1iXb/JlZptsn7mu+LV6VUp3kQj
caKVsrK8tnsK0kt6MGSqR7YsUNcrmlSDPTOfVGmUIDhH2y42VhgGEO6mNiw6er/K6SQmVNKGHHdB
M3Fi9baBbrcr1YhqawL+Wp9gfuTba+LUMYUxczevHF9vadVMsNZJe82vrMr9CuvH4q9wLeev/0wQ
LPb5dhYvQ0tqUCTy40/vI0vRc54jvwN6/z0QFsF0mSoulr6//YlT72InbiYapA20aA5L5c9SnSkj
tTUQ7MR5GZzgz9haIxWBn0C53TBHfgs2rgS1tl6PNsjDwszHRq61qepQGZIqfLlKh763dZgbdLcp
KAOtRKPhWYrc5A6MNViWsKUlvI/akr1tsEb7uSJ+eC4gRZylSZzBEYI6hndOu7dEKQOqga7AmZrr
C7fUm+IaX+YJOxqHNPWPKaukpEW3syjaeeE8paUtIdY+nksoUl9kYljrPqd+XcgmGTeVy+Hx7nHH
rpB0K46dMVrV5CEi0tasWW6JHfd6RwjNPGrQTP/enCNvsh23r3FpZgRDsYQJcLn983ihgVR8PHcF
KF2w8cpD0vENL6KWkDUxRSsm+2ChfeGPFDCnhtkCn9Hqv+6P60It0SEAbbxBDoJ91Aj+XFnr8XZv
Zf5ogyEokQuzxOUgpGDM75jDiiEOik/K/jO1kMx+yluY9JlT+85VU6TqpDlMovAY+woEIUxTUHpW
jJ+Dy0+dcNMzuS927tFEi1d4Hp/s/FFUI00cV3RR+OHITYApZooozDutXg2hcHULYt0hgI7A8jQ/
eDwUs42PWTZXIZTBB3tYcnG5yA3OAL8lrTgVah556+9iUGk27Mtn98cUn9tZIaRGVR1T/lY/naNs
uDFHD0mAHhVlMVshxfWL8R9aGoK817/enq/WnmE/AbmOUXihs0Wmqia1bbnZbSd5wXryoEIaIFRq
xPnGF2IxieuYZ31BLXEbr/2KclmP5bDS0boNm09z4h89PE/8OdLxnulSSBLmqYXBMFhWRzzMy+7Z
qZwCrLBce31QI7tLoTnDoa4U00bzN/2Tqd7/vtCx9czR39UhTrL3SzSuZ9iLYZHduyZ+kLEVztnz
o25eIgDP6Pt2I4s7mxoToMHnrJZUYcryNmk6LoXgMh6ePV+oPg02qmtVyFXZWBp+I5wUk3wpa3VI
IugSTm4aceyuk/fkZRjcrsCbyptACQYC6Z4iZr1aHNQIA3vA9L2dKtHIk2Fg7dETBwUR9hQzP7ow
rk9izgHXUpdZlJEff28fChj2GqbBsQVtO6igCmbHLW7GjE+555Bp5SlwMQ2HvTjKAnoB12odHmPH
1hNzBIcugYfVjASTWCnwJpfHpMoO3AJu5gLAUBEw9d2KqCKCT7H8JxRwUxvdv2lbbeHMuMrkMntD
VfvkOPl2aFYDCnJvmu8f+7riiqk9q2E0KvCQ9TskcWO12SWAOrom2QN8XJ/CCnD06NCtsaarHSba
zI1tTKqDS7CXDtmPkU1gbJngqgmMN/mYRCarRFqXm+Mea+zdAzJxtjhKmu2U7+o77FyPmb8XhRMF
ZGE7lLELLFRFVbBthi0kLSRYnpZuhqSspWQsE5nEu6PAQGmGOiBIkEphlw7queB5qn6+Hm/BTPoT
W1IdA84eBO/bXSjun88so/8UWaczDSEH9sWYtrLjf7AEGRTXGQfked4AWkitpoJaXVW+CCG6zeXS
DyF+QzlcS01UBcfjckggnIPxz1KfDIFK4KIRRAWfyTVz80lB0GovELX90U7elhFFSXpWZsmUAB8C
ivMtKRRkz2sCUcaGXCEk0oyKtgPfEXvRb6PjfyhYnKTpeYfH447+SEUDXzRuQjJWgFmJLjWuTAkK
aKRpSA9U5Onrk6hya3yZev0w2zS/ICYOREdonykly45N6+m7+3OCGH+2gcZkOE6OjIHRPIKO14vf
3dnU1Wwe7PsvImbt6nUsQk8rmq4FBYOBIP45EVVizEZS12gHyo8HkfGXDfOCtKs3yw5yqoxL/Zvz
WQOydI9qM0Dq6C/MdDV8F77TVYGbKGKUAfBbDk7pCi/NIjNmCXK2hQ3HE6IqgWY+5/YA7YV0vXnF
XJhD5h5U+wruQEbYlpjImG5wPxV/PyEAsozU+HasR0QcgOnWtXvGWDHG9DJYh23xDcsTE2y7etl4
nKJJ0LQ9Sc1UBDAFtCJee+QYItQgpZ/raQy5Tr6KkvVzLG+q/B8irzHnpnQZJL1be/GxoSMN1V7g
4+LfHvwKwsfsCZOn5qTmI9jHpfVrJzRkXhuJ7ELUlZQVQ4YU+P0ZWTb41922PeMLe7Evi+zu6RGH
YnAQiW44q/QVvvWGD6PO9JVI7V2Mzsv2FW7kxs9LILT0njR9Fr+V7cFOZmPkHLp3IaCpgIrkkUPH
I/qAoDSgH6rEBTLo8UwndCMawuG+dMELbrqp3QhpLP7Qr0PYjsub15IbOtAHH0UOvx2LlMaL1Uzu
KzTQc8J4WFXRe1UD+QfVIjXc7aQ3J74QbMBjQY+dZSsn56LWeGZOI1d34RT1LmUMon5MhzJMFoR2
vvpH2qNZ/P4e620+Vpc8qqDowTZTtXwon96YY+f9YdOi7ShOw/5bo9L32+CepW7sSqe5nTn0Emoj
CvHk4rNBJKWcjWhY+Fp77NJFNxyhAoxbAhuSJIsxW1GCKQ3Q4Mo3NEWm4JDFBh9Jisv0/5z7QFQY
mu7F4ampBYWPJha1E30/Bauy6DQ8kfZJeTtn9SGYdWcTwdkhqR+Rkn4h6qwhrbCC8Gcu1xR3rhhC
8ldvhI31QdZI0PjYni9cMt4BqM1/gf3sFggriUC1Neg61v7o3RxQS7cbLUXXdOJb54Ngk9ar8Ipo
rNB9hhyp0m+OLWvQe+ingxlh5s9CVyStP5Emd/yMAeBdKaPG7mf7tqComYQw+vmQwBeosLNzIv4v
cTwd2m8MyMJc0swbcJ+skwWO02hbBQIgEuT4eRt/rIoM+CSbdjtsGZHtlt+UPJICriK8jW1W6fks
E9YXlHSA7A8kXjoiqXBfuplOceLUSSb9/V5xcKkgNOTNY1U3KPGXOE27NDLo8iW9LmqwkbcjxJ5G
14dnQiRh+IUbhvVD3pKLPM2N2XjS4y9tDKLuAzQ/6T49h98E9OSknlF6dAARwJ/EPPp7EGA56s+g
M50P44a0NR71jOrHu7uob0DfjyhMTUXsY0vcDIZyCsU/yNy9znmB7M+eV6pmtYhn18CxaH5XTXVL
9PkvcvltmXoHZ21z/n8pUDmU4xmuoqonI0gJrKzYU0bWayPdGDzXFvvu4FzuibpG2xdGoC4OIn0R
wHmItFdZrVjAH4vx8ddrFgvCJNWYbats7UzZsTsuArusVAgjYR1/y5ycNHhKwPKoo8PbwNtFIUHZ
dk+CtL6hlirejuncQCBjKcj3B4MFABrvgVHV5/sjequfX5GLDar9zIV3smXVCCMjk70ES00zYs6Q
t2x3UhzjnJz8Mk0vi2H3CRuw5Pk634E2QjzPw6HVgIg/0rOGY7C90ojar8bKmYc3tyZDdC6bzya5
+fwIgC6nls8tzjbk9WdtsgpfHFw7seHfwbRBxR+CIVSO3OHbvyAnIuf4wag6W/KrMnexpmqscXC0
NeKecYyiBaVqq8IyHHztRelznbEe25X5GCNDSBQYLrKzFbITtIK1LUguWsxXhKxj8tPrRXlzYjb/
VLumAn/t3o6NpIr79u1/fpd9luTSXi0EYkpRzNPJzf47aKxfk7SvZaPOK2nnzMy5S6TmLDBCuqC2
JWKPE1wzFdNLGlInbzyiudIhCuj5AtcEZE0rBEfCltdoio++bnUd2VrpM3dDbu7KJJmIyPDtwzOe
XFIGUQeSfYrCOpg7Tta830by8l2CLaUze5tZvqSx0i8LYe+c/HBsJGWfxI6Erc9dDzzXxB5sW4WK
QixADjAURMEoqHy00GlsWlGPz0dEVK1PJfYQXokyOS/nkfc9wfKtAuGd/pRx52Bf/oI2AHp/QlW9
sxYBtO5VcdltLnSldG7fQM8zjFd6AMmhVMYQ+daxVU3+DAKhRIriJq1t/c4/fl7V7udKLzPMPpkC
uMdlKYUQfYfifKHGx7O/0LarILOVbT4x85VntUSvi2s8SbotJmmAxoPqk+8vwX88/yILUJsd+NcJ
812dsddYvzswlJfknNzyxKaMyP74hPOlUO8vCreSvqIe6FP0ZknDGawf7EsNHrrkyFIfHxo04dQK
pfqXqxc/lnqMLpGxOs2+M+EULWpcARPp3ElMrdeFtX3o9R6HCmJ4yI+Y0sUaXr3ajU+lDPsFskLY
fvfw+gu5+gmq4AvV0sCzkrT4yDBPsv7QdmrLzyaTwkg7v9NYK+eQpoj4KZfxrMFezdDwsetb4P8V
Kf723/KpL+pAdR9vE3F6kVDdXAoQhNVlW5bcfmuZwifN1JpVEeCPzG0/wAp5DIi7bcR6EjeQR8DA
uU46MGiEKC/r3Y9KEwLZfqED+yiW0+Y+dDGraa5VpqFpTiNzaKOfPTHKvaHdUrXTe4H6GZZ2TocH
HEED1/ChhJehQESEZqWqKMt+eCLDI4VJhn2F14cwvVU8eORyslbqFvaNO4L2M5LtIMusg8b6HPhm
xkdCmyvQnb9JdDIMZ/K0Yu3HevnhrDrvsFyrSFzXgtVjrUESWWt7T7DtukTsFc1vtsvMGnHyrEyU
FmpyMO27uigtY434261snbhmGIuVUEI17fij19zMms1xmEnaJ45eJYS3k+JangrWobbxb8dp0bhp
3KhdUsquIhfTkbjxaktOpACh1Qw8/Lsk+TWyiYWGmcbrY2vpnHidNsT1V8X5k8VRX68s1Tvi5/iF
8txmc8+J7xtfzYqijrHcoTzzCsyHnpa2ZsSByg5+xRm6qMq1UdorW7yGRVyp65DOGGIBhS59nc9f
SvvDRssj8GbSbmrQQ3Qp1Wa6AKbEu4mYMkl2w5un+5HLGOUTl4PDpSnI+jgIKyWChQ7QFtZUeGCJ
DedsryDzbYQMulVWHbbeE01zJUNnR3BObj62AjB9gAqNobICFD2BfM4HznwziVSTO4GGXsr8xko7
85aTApU1uKt4V0S7PUQPE/KKuexvKaeTIkdv3zjO3Av3vCs7fbwpZ/Bhts94s/bhGiKngj8fk6st
4rglg4CEa+3UpbwiwaXqjsCoVa+4D16zLfzkF5WGwCrEwz0nMhd43mHzRQDwt0SeYytxobJO+a7h
UfpljGJtHbkmIh4b2Ya/nJLz5TittUAdhBsIuBbY2Welzr+nxmjR2WDhVpU3nM7zJO7KftL+k7x+
vf1Jgzgc8WtAIS6C7xFjJTrYV4Y7buF/mJdS8DgCMB43TvZjshai8phKQgOguktvgbh0nDtn5wsV
gFJRAAI1l1R9MjnPweMQSFIpkFsL12758/N4uV1jva5dCRtkRNdgs2zr37WPcewQVK8zqxW8o33O
orMVpm4PO3uN+ibqOVca0jQ79dmrrJ0Dcwa5so5bvIUQWfixZ2dlzEVg3vwJANFn+nsqvsTqvJ7Z
IJWiIFF6JEQ+x3N0TZ8q8hi10hhYHMsKMK5cVbwRRpbqF8P4REpqTkP8eBaxp+0kb2dUzNFvsqNk
x+dwDnq+8lL/x/RW8M8odGLcTAxz2RJcKyuYJykhYdqhSnUckA9LrAvfwB9Zu8r6rm5txH+X86+o
JtUAxQ3WsdSuPaWNVTePplbBRXNut8iKWn/zR0/8fkJP/dFSC/iQ27bLX7jAGx9m+5GY4Tdn8gx2
vVLHUTXxJKY4oC6Rbd+Fs3zM8ywT4EO6/XN2sIU2TkAMY5xWb4pJVbajkEDY4AznLN3x9lomJdBP
iSLj9WsN6nbatO+Xsj8MxZ2EcbGus9rMtcdRN88BxS2NqTvMs0rpGbAH2NoBbyuYat+/YKwBiZyG
exazxuOWTprR6eUANO0OdmeSvEAKjMoDoi0xzYxwMfayjmNmK8qaRjz6QWaAjrpUppqMwDhfO83P
HgggLEKe9Hf84bTQwRpQfefMqaHusV3WNhbV5buphEJj3W6S6TJXcEDj4IkxvWEsx8GZd4pSug4U
qWh9tnyN+617ZMBxU4vHhrddhWYNVJM6cpc+yWTQEeNv26I5OnqYh5bRmmOhKOX5OEJjnM9xlbq4
KH3B80cHujTqd4GYn2PZ6Qr0u7NwVhYzr0/GwvlwKPURqTY8zcLGZ1nyjknNTtcHZ77/chMEsZ44
Kfjl6awn1gX3boofQwDx9dWwHwS/kM9YUd5OEnXKqoRBFOt9TsEiaN/G0gKtowub4GM+P1h0skBe
ClJGmayI+rDkxqhwoA9bdNozPVu8bbxtgnQEM7ZrWsX2qWpnESd5SEYsHjUTsM9Ny6x3R1gxLvEv
9ALx3JzGjPNP9vb++rqajm07bAi+1NWzQF/U6Bj1yQn28ebh62DicxFeLnz2Tisk7ZwZ+tIpC86Q
2MbnaaTOw+2mQ0+HtZ6aHWqrb4Hrm07IHTAw5dauYv1ri8ff5dGcFVaEuWF5LlR4GqBVy5cuJrc4
6f7mUFGKj0E0fXXDN0iKiq2Dlrn4sVXJTVaRUuyluiWheTdsYT+oqtY2hWhWWy4FuOU5bRpwYXqO
oEzLuE6HOwSRQxNLBepPPFKPfp3vu75OIG5e9xVOzEQKBHBPB910btVR/N9//2PNi/bBb0NluiRb
6yG08NcZkhcyWHM/Jwsb16eUkiQusjqhMecRb1ZU0Vhwxxx2TNpY8Ob+JiZhrytasfC3pIQHRvrV
CZ3QyrVEtdHYDyGHIcY07zSSbPawJ22CzrHYWgEh2Y9Gy0QD+lCUmHpdZVhu3LQvO/tDhPTm60xW
DXbtNhxg55ZgibcnOerRU2QZxBKLIbbs4WvZmr3xOYp+wkGhVlZ97YV52WGfJ63iB5lnow6jdKD7
rt8cDwuXi0qKUJtvzYa9Wfymgc6W3q5N8o7jWO9UUafomK/ERReerJck4vvC8i4Ogiz1JVGztkdT
eIuV2EgruN/1YiBofN74WVIcVMx9xwGKptfkrDX/wqncakoXrGNTQQ3xamSGFcD3SEfr/g8qHA1l
Lw92r9VsNtZaq0wM6mkdx0MlcWPVfQBTCQAOSyZzhTzsoFWiHsbGKQAztkE2DhS782QlhBKTtGDz
hWr7NJnHV0WbfSknJFvnas7YceqKR3v4CDfe8+w1sEZ/rHriHNnzAh2hjf3iSXprt78m+WEKRjU4
8Ge5RPQP6m77v4y4ggDZ5CX44Ysk6PvHavWAxH/IHLDsQSUVKwHz41jWypSJ/y0wGXEczBE7Nm6Y
4enIvoUcbGUD4kafDyEF2/c5G9FXH/P63cjJlduCvazr7sih+HizAHJDTbYPiHGLfPD42KblLVnv
pH4KZ1vH3iHG5lXnHckRVfASY8pGyrrC4drPvPu6dw0Qm7/FIw921XmNW4BPA7n9ZkP+dFEuLQiP
cBlcA8bl2g71SihFXriIGoqpKDouDDg1irF+dKYYIuvZsMUNuybRcm9/tlmDuSmAs7eMm4cx7BoZ
p2y0tp+1GuUmXJsWHXQ9f+4dJY3ggCr5kvjk3QTjIGrjvBcKJIUzIrIUqj5g0WVdKj+J07w6wtf4
ZS7btlnSKAqmSDxOuGIL7Amulb8nu0xqLIflkktC2gY0NxLZzvpVAFVWABCLr+vDHhO/PEQAApLR
sFbVMn+bd0AVsTQUOjGvP0Xe7ejuShYKzyVjpFQzQpKj1mYsRIrejeGC+D+veMADjQ8yPkmNFC60
5ij2df/Xkwaq55HbvicvLd569ds3oHE5iWkHKyat950b1qYQ2apONsBwZ5ocHApbXZerr7FlLV3x
A+AMJ64gnmAAKWd9IrM1AxZHMhbw24WcVirIorIcr27nVeJqwRy/TVG9TNGPEI0G4xyvUmgvJQ3K
I5aJrXKF5ObkzVy0w3mFza8nnyjHckF4NEsQe4Zjhm5UBY24FAJmNznhbOdIOWPZhtobs+xHNFky
Q1cBy0pvC+Rs5jOkoP4QeWx1iTLacRDLeinU0OqdcCbbpl7fFB3sGP8NbAMV7wWj+WSgbAgImfuz
G+lGMT4MG2yzuHNRsfRL0CLX6i4yQ9li5Z+ou+xiLLBTl+6fJN9zuFn89ZIMu2dZrewl61E+uFfn
vwi0Rc7oXSccF6AYgCskJN+oU+BG8QDCedSBCItwZQvGWf0wAOxVqw4iLRAPc2IY6UGdQaJfQDDi
Xk+VpWUNCpkMmD8oVXgNjwPHEM7JhwuFfstei8+jbnQYxEYV/J4HwPXKL7uOduV0hvGumiK4UNFu
eujcyeOnMG/ELjIuGEkteREjcIKsVz/vY55J7+vzwGw5j+333RUaOf/t8Zb+xZu++DdfdYNuABLv
uugas08XkiVVfOlDwr0obstLQiwaI5+CcVO6bP7bf5Rudo+yP8BFrr933hWyY2sU+WobhHx3Nxjb
eRpn5VSnmGkuHcp/mtyTs07NaBdFjHe75sJtpEH/Oj2nrklUoT48VPejnDljFixV23gueXJcUAvE
ZMTBAdxp4liEssTQRurxXNR3QdJ3JUztUL0qe2OdEJe2rDmF3fWLsyUrwxKjqIXVG1rMkPugriXt
nrZIFur+eHKq4EWWPFxmCoB2BLayb15KS5fcHHYq3Y4U7RTcWtoANHqAbpOpLUeX8Egjm2wYsoDI
aFrxhng2gB03rB6c4DSSpnprwLFoWj3sbv8ojOOEk56GxgvxlDhp5zBlENighmtHN3PgDL1IZl3s
or7VWJ/XO4KwghVMI2hZ6Yx0SRRpVl3EAT3EXUH6l5QXX21fO2fyvQ3c4dfjA3WUUva+n2Me/n9p
klsR1tK384kDaAnnDO7m3Xiy9RkqGKvJ1IZK3KC4X0adQwU31AxyCp3RGskfFX07iQ3TYW+uXmtZ
Cxzxgd5zG2XNtqtuJYzSc1bAoMPDo8WqgPpblxuYXE8FwetxQcd4kEgXHTMqpjDsbNKQPQSu4LAU
ATlFsPF0FZ4Tld5v3gqhhtjkbQg+0hH0glUP5mrvfTpnzXAHtjrhyvTapFBzdchFjgTA7yOIhmlP
9geJy3PBepsK1Hj0NDn8H4/h+qUKsw4d8wEGBl+hORm6mlbtCI0E6UlOAHmpf/Yl9lZzxqZ7PszH
ea0u+AwdZ23czoYTLbY1aXHB6GLj6F1VdPNLldZ279H98shtJF+0DOcQVTsxzBoSvkRfABw9BOg7
N/cadi94mtU8Fg1GrSD3mCpHssqtwTc2jrtDsQrdxMZ693Bur7kcKByZoGrwJT1l5d3RKEb+7ffJ
iaLhJS8eOkIz67nSZzJgQ4Gj6ziWRVFGvpGrMDifv3JoIXRFid/ACEv6FzRvRpeaeLkCS3ueJWbu
t6ZkYVw46ytuGMrGy3QDHK5dOB0x7yEo3Z6U0VvOI66JFB1UfYebbUtxv57fHcdF9evSB7JQmpX4
sHcCm33aHbC0QLc/UhSnto03CvT7to3jL6G/05B5QPs/dkomQ0UEOI+nodAPq6UdXr6NZuotst98
XBNbU6rgmcac/vOaTb9+byQ/pWlHWDy858tORkzGlaPj6ScBvIONEQ/PxGFqHVbOKFx7KQBU+yMJ
GZBqwLT2Gt3Lqtw1cWFZUfa3GtL7Z5nwzU0vINMa9eBz302D/txen7mXcRz4YDTVrFCdCAcvKVzd
snrVw/xco/ZqwyGL8L0/ljzOnuwk1gRIL3RVZ0T+DZjJ2KYcar6SY9kbOzV4yBSEprdywHJlAbL2
/wOHxm8+h6lbFT0igd681vm13DlWVIIHF6BsUQEouDtq2uWtzjAHfjiBg8pPjNx6pqxwibbycolW
EaAPw+kqq8V+lc8gyN7CiEiX2DIX1N41p2sHHsXlH+uGYgzo/J77Kus+MW1x4vZVCsnyRLSEdLN1
6y34ubSNURYmRLfYXxTwalGGKNTKCpBo39XTyKUtoJvaFO6krYIOkljOyOZbEflRwNJfAJ+PFbRo
cIScOJGCZ9Zv6+b32y9hvBQqGEXwxCzTr2ZeFye5HxPTm2PcTfaGusWuVZIcglqHw/NF7y/w3EeG
+McbBrfGLlRIUfVPrCt8Iyt3/ZOOgEYDabsdjp2PyQzez3es6AEEsSx3SzLm3sr0iRjHXWYQ3Aqd
weGXNvF16jLkHgOinsZ3Oyc+VM/dsgVNypY3z5w+rc+aSxrD/oKZCdLDW/k+seHK/wIOsFZvaRJT
JRY9P4GxSjrS7bpka+dDlE4hKYY1OhWKTigbJtMRNUkhRKdPJPg9RavTKkBer4tT6fSlpRiPUi7x
kbaWzylpy8BLAVXGnpWbAAf6wsSiv5YFxGXVkSUK93QLsME4dZ6AfbjJXmCUwjsjzrcogmeitEOB
bU+nKShXyJkNaslaP64Va/IfEKEFq3Rk9LdfTgy91aYo90iYaMp8lYpJOaAnY3gcfMtsGbAlt292
DbnhvcFYncg/JND44E4fFThRkcoLUc391lDnORidgJhLEmQmxSyyvK2YOXnV69tYk/3UlJjy0ZbN
0VqL9NdCNMA7jT7obduQpGDaUruBUbGPJVtLVuXd64njnLIcnRmVf2eQb5nlNVgSXxurCMyTKKsr
Vznxt5NsWDkC86DU+fiI2/iJ/6NrrS66+ho4m5XdicNZl/NB6eMgDMZ/6YhHLZpQzr6j7bIKQpqm
H0BU3keSDjA4d+DitUsJHVwJFkRZg1nbCMy4pQO/zMLZ4Sfinj4L/HEx+fpkjtRy7UjwAjHIlWGK
uULN7teXfc7T5jcUZsvCE7f2FQbj7kZjqr3RIrkmknOOH+rtlxX+il9tvzx0bcpL3+aR/hmx7/bf
K07E0Trskl5SX14Jq2W/cV2RusHPdTlLP+Yj8cZ1wghAVxRFUNWvO3UZWdCL70FI561E8fht3YzF
TA0Kvm85kqIbxoIKiAY3oMHjQdiiYxrZfBpkBxjTb4NPNn6AGeccC77DAc6SCkzzS/Lb0Arn6Oa6
ntDsrTIJNes4nl44mXbiIqws8wJyEEjrv2ogZcCZBhpIyTFvRbxE3L2L8wZpj9LUfXdI4QopH60o
igG75f9snPbKP+1IMrN3QDqSJv1YMrCDnLmRLDblvAqFjUvl1G0s+ou9H2BEpuj3SF8SiR55qsI1
k6i3lM/CV+Zdvxmx9TWmhpfCOTeXYUGPn+YY97nKDvJ3erSYZ7DyEaxvPROP8NHWEbxlFPYBORmp
wKRnCORkeH40kGU/BZ7WpfEJqcGE2MNGJK9dI/Yx+k248WC+nOvPi2Ozh8XtNnXq8g5jdOxJq3C1
aGmL+1nG7gFsqePt0K57xSPc4BXZjWrr1pxQW0ZccrKYpArz9lgOS7nfWOoDvhJ8ExyNce0XnoS6
YSMO5JWQ/bsvON/xXDf9wgSQ3R0Cyj+OhnUizUJU5vVgNsTP8NjTUxl65uF1DcBOjJLaLgSnSA/I
woW6yNiYeH/3mPY1QLtKY0RHWML3XoQBO10L7pYX8gMhqfsnJz4qoTtTDI+cP5RoWClz8ljFegex
N8V2worqff+C+xr0PQxwfkZH1FllTMyhABp9XiffLSW6k3EVSSMhDFSQIeDXVYQb2MTZBBnpJRKh
jY3j4/eSPIVAsrfBtGyOlfIOuQuRlhHtRpzm2slaLsMOTVnhzrgNQGIKEOTCIYIZK3spyJtrdEyU
rXwMPRo7zmR6FNHRNxkGR7J6VAKhW9ImEcGuGzUTXHZEBltpoNB30z//AK7DNG550t1WqYLHAx8Y
kwipveaTzntWja5m1zHZE8qOlUmELs7B6FxykbMHUsD687MAILTY5Xk/cNLSDrCkxNpzVfdUOd34
DV9GK/yv8Bgzkb029wIfgvu8VakyAlwlLKrQf+RbtuVVcbbDcDML+FIDo2Nx7ryMX4iYqIQ0YOoL
ro2X21xRQlif/63QZV84GbyFgSW1zpjP9u6pQB0eXDbp8IB9lypXIS1qxLfoCakWkIfHovmA2i1D
H+kCdYUMFsppm6DbtZDai21FQYB/4+XQtm14vaezJAf5oCdUkSggR0IUnrHSUTlFLU7e+9lEoM1p
jfnnU1Kjs1mjnSQCpU9xxmCZBar5RuJpLY0FeQeDRIs1+4QeXYvLnSsK3pL3GpyqBFz4rx/xdD3V
ZRAchsbAv7sB4alVqO3VhisL5iLcoYwG18VuUE8SpUNPt/NUcesv7dn0RfwzCrFUzUSUa+eFnSEa
Tuxeyf6hYezMR8zIzObHnZFhQNiTzEGkYWMHeB28WD9BaqsClX1QdWeynHD7LDw8dPjgXfKIPdKb
imUwtDDTVnWWOfXDmjOi0pkEwDn3Ks3BQPRFTAFkWHxQ20krJT5n63qf0eJ7oXnIgtGFqYNfKZEd
LNZKlnc5AkpAxbSv/jJd/tWxJYL6JBw81iofRbJMujS4eVOf/E7PUvx6lWROmXOOu0MboqjwSDWN
Ya2CMF+53IWTGtgENVCA0Ed5+dfzXVUAtAAteNeSQZlTbZZpvu726UnEcEU3ah1xCOail0AcIIjs
nb8Ew2h60quZURTUKJ4TLk7a8RbQYcvzyusxwCx8I4/ruZurfmRBn5At/5c7i10+sahB6k5uR/se
ONjsqxsM7tJsjgQDF7jaiBM64rKx+y2iCTAcFCDovM32vWbxQnziaZK9f1LC4HJ3JlCR51aZh8xH
ObGtf6gY0Rjd7jwgjYpmC4fQEuql+068uqPMltLk0E1PsvEo3TlQTB5QabRW9jkkyY5/tSsaYy0D
IWR2zeROyhtahP6xPsvU+h0kvCCf8jrFOvglvMXjfFkTIQYfxZeRTfhY6zs9cWA391ypeNo65vGO
caR1/H8VIum2tOqJ+Hfx+vGJEclbngyYp7UeBCDU5PCMrX4V5p3M8UZqFkSdSl/J+ydEDOU3tdL4
NbahtJC0O6u1LPvTFoJZDzpIiO8FRVb2S2G7yS7FzIS1rjn8xgHWitbaYUv6TiZvbRxUT0EWGu05
0AxrFnQVrUlWTIjtYKxAvzsmC+TAE/4Az1h0KmiKjOT35KbqjtLx1pwLde31f6rJ+F72BLTvPKKm
rBbnhTy/JltKD2jvvUWxGUAaExGz8/1pP44WPnDuAABXhxMk0rp/spDitxajbjHwaIFBK6ly3m0A
fubjTT0vfhueUpiDOFHBTbgmENbIOgiafu+BuEjP5Gt+i4Zau5rLw+UB0rdFoMMAYnBy/C0zlufh
hkrSe2t8cdhZQub6Pfp7XN4vtol7+S/OoVJXw2Ex4jpvTo+W0eqLtAHIMnaQiEgAO1UTma7EMZjj
FJgg9I1BKZvGDOhT8H2Hi1/qL7yRt3BOq4NnO4G9O65p5q1T1vpbCYju2eG5Bi2gkifNqUScbK1n
RNYp/0YMa7cxXM5rshnahvlYQanRixkbeq9cbLHyP/QR34r6HkWWj2LQn0oNAdpxYrFgLUi65g3s
KkaHKb6K5AZRLsH8cO1CsMUOoWkg07lAGkUg1wRMYBd+FvDagKpgm06F1Pno9wW0KwXsAvOpJqvD
Hm4ILNygwOyob4Zz5evUvGAYRUBEReWFaAkJTQAoCzId6XV+705c49ACiHcA6xNYMuAfwqVnbF8M
zsIDWwjDEzaC/Lt9Ob7lMyVgnMotrdOyMvs7v72tP09MjxLpHIBLGLG6cdoQSGXfQpQHc2OkV1mp
oP2f1fSDjoFDcsYsupoF7uaRD8VYTKbaYOjxFgKoYJl+TQHQ3Y+7yxf2rYLF/+SZJRwimecmkj5f
HoMrc2vn4ihyMrUt6Fd7vqYzVr0yzMoYv2CBrH0shQTBtibj65dGySdSwjg7hX2slnheXLCqu9yT
Mg6jbPpL6TX1gi0ZdiCCr9U0AR8gTmohh2h4Ty7h0NTcJ/hpU6XH8Q7nWTvdpU7cHChTmYg+ut50
Fl2ZGOxibfCkFkjsojUm90sYIoicgd5soI4pbvMRHpxaqj0stw/vUoatvpsRPPS9106JVg8Z/IBQ
tLg328pjAKCckVufgkrBgqVa4gt3IPAVybAN8HKEhIERGPnbLh6YNVfmWUTw5QRdsNyuPGmP9B6X
MGxxaVdMiLuzUJLzE4SGJ7D9lNlOBx8nDYbbsHpvG68csMdv9OSbddrT1c2uNx3BXkU9HsaOYgeS
fzeThJfFSNilYMU/XzVPzh1v95LnZYT6ReU6YziJX7H1yD3jc7Qqfaq/JViIpNJCNp9pwo7DZMrR
psOljwDnYQenW3qvFsQYYFHdquwokDByNhROmHaz4MiM71Wq3O9FQuxrdtLiK88bXlzt2Q5aEWJE
8XWrbDdjkP7ujFyyXsGXly9b4FGIcwd2srHrgcm0oV0glBnpTrfDjKdPNRkzPEIzA4NGM0K84TAW
s81Rwv/dD5irF2dO2jhPsTYDAmyImEgZyxTJiExr3ML9A/nBJnq1cN122ZzE3IBp+gEAAkZvgZpt
8CbbkvEl60ejDSxii8vXR7782ibzCHDj+PDeTuj3YA0iw1a5QRSdKcvaqb19qjAwtz9dA4z9uj7w
QsQctJDEcuiZ29+UXO2ziwkescelZo55BeQAgj7zDNab0vn3Qc5Ac2GyH3Qmj6aNkmbYalAsHS2K
VNYvAPaZq25ouw0xsUNXyZMelGIPgX3qVdSak38a8ZS3gtFePri/CMgZzcZbYCdvrvEN/NnWrn7q
LfhQB4mgXTkkr17JwpXmSF5f2g+3o0/0H9ZXpJCQxDRj6JB5R3lZEKTltZPYH/HOsaLyYaPNsERn
JGh0xW+0T2PK7GWpXstACY73EZeOwWYRb+/ZXYbrabSfg+w2ctJq5LQCV+9eQM24+RnSNg7hS89K
8hl3eESZFA346bM+t9IFarNlliwL2ofxZ/y/bPfs9rD0icpHkKUDBtwhiBhUVnQpDhXd+smToNtm
MPgHjFmxaDVD+aBVp5AyK9A7UdMmWGQ2/j793XqefXfRuaXW8nFk+N+xhws3LRsVd2qEKk7Biy1D
CYQekzWQ05y3oquVVmFKdW1SMoWAV8P3Yzi1l3kpLFq09Rn+TRyKQgFg3KxzleVH11RFHnrbR/ic
JXZhox3zubTPgcA/AEU2pR4Vfuh8VsuykxF4J7FQC9Hs7lyAm0HTe0ZX2N52IuHf5KEp+TBwIaGr
HYd06s7Z1wIoX8HMz/C8bMm9730793D9P1iuB3LSeKGzo7eZVxLyrF5HvN0x1dGwFTfyyj8Ukv6Y
5M0sAKlcUrI+laNPiH+8o/KacbiFQCeNM7b87o2k0im3Qg/wlQESyKk4TEyxNvHBC6HBkc8tvObP
xX+z9C55vrTc/AxP84i+pB9kuJvnTnhedktiGF8wnGqZC/NJ5AoD5/rfMcZAnlzn+15XTrfhzrgP
/ZcjCfT8PIqnGlNuokGL4nPpC9gJshdm12NgeLyYsz2WdQ7MaFgEmTybHmmb7eVXkGEcNiDNDwAS
kp7eCSu9Hw6oWPYQlM/gmVsh3QRNo7OUs1NzclNEhU+TcsJRh77V4A+qA7y7/sTzrTRYQU3UVvMg
Ok0NGq0+G5XUPJfOZA8BCbkzGuOhJwKwyqM7xPfmC39jKD3zBqCfkU2vz40/aQ56M3CIrgAb3cK8
vx06D3o1pX2mC31jnVhjq+56BcqlGOZwHyjx+4/gw4YEk9H2wuut4e9kEZBN80RG4++8Fyama0kL
VUWyr/lV/8Q7ylPWHoKNg5WkkEd4kIEdMR1/HPsCP95B1Jn5EV92GslyOcSbGdQDGKmun2PfRJHi
hU4YwqTspfDOktQtzU7yqED/J+J1vV8bOgTQPhuwWuAC34UVf2XM63F9mBCTGYw9Z8rga351O9oM
wigkVwoa85YEaPnp1lI8EDoT7N2vcl/GKtJXU9eBBRIVU4KRlj+jlEJHAjROAJV3IxYt3XsOi3nF
QeMsRMHB5h8k5k9HqDN/aiRn0TDLyDkXK3kSOL4bzn+Ie6W8GRsNqy0GG+Rx0pH1SFsTPdr3qeQM
/7R3QzntapzOhaELg/bDqBUaUuFJYsYLjikhDnYKSp/j+bEwFnhCiyJ7ndOJxrROZrDrL1lyS1I5
Qlg6rcuD/DJeuVcOb1JGDCkykjGbZqAPcd/Edo2BpXlA4+tGimcGuFbM1mkSlCHlRBdEi49/lbMv
9I1FxWLfrvJy1BUC/yc21jtVyI65sKNJ1W1LM/qJ7ZxbNVrPr3WnHL1vc7nT8eq7Xfqh5r6d6X8C
0CfuY2mKYwtGhQoL7K+GCxWAQiutUIIQJcSX8+WNoaa/fd3+6wZ19JBTn9083PP4jMDDoVAdoAjX
KQSnD4s0jomZTVLej24fvedqGv5vG1d86Nu3kPB2haQCXNAl+UKwqCDnFwv5yBbrje3QHQi4QeWO
fsPUFGGb2An16akF/QMDCSJZv2P8djorn7YLYkWU/2zDj2Sfra6qp2WXFkj7ut5Q32uw2n4yryjU
l+YKSjRmMm7wsCTlBg2ZTgin3Rhbiw4/MoNd168HAlCFOd/+CEY5l+7jE2FbppA6Dd2oGMUHGXz8
ZRzx9tOwLTMZVoWzf2Tsl4qyQkWY66XW2MthI8vp3F2OnU4mOtTsISZt1N7alQLb/qfo7rxusjhJ
g/KMHFU4d0KlFRuX3CkXOCCCt7dMw2/I5fDTkDYkFKkjOkHKTW9Xxbkk71p7ioBNQr788k1wx4k1
4ZFNja1uBKClZbEMmgvCHWHBCmHnuNEze7pPqPkDyZbCSSVXzr65rBvPCKbASbrEAHBPqw7IBVz9
MTEWeUKSbmHUet3pwchEXiZuaZ3oN3g0/0zik8KOy54TIwFGc2xZvDUluC38WAvnQwj75rgTzBZ4
oHxnpglcQU/cUMAPH2fADw4VJYavzplba/qGtoS2HoBdbhKbveDQl6SkTfNXm4eo9Z1HB7CryVfh
hlzvoLqcsa6sZminqoe+ZhZsaYL6WOa17/yEee35+egHcGtVvVIMQ5fTArk3PDZPYNKwBT8FDGx8
wAVp+kPbVxUc4e2JhOMw+46qZ0pB0+xoe9Gk8+lX5ZcU1Kmg1NY6EvrMOdAq/kl6BYDDoCwyTOy8
utA4523vHA2wyCn2Zvvxez9IUb9NcIs/dJ8lQ1lFheJFAjcNk7gsURCioadLFkPHkEU7jbtbC6xW
OUhtEXCS4Rra84725QxnVx/Hvs+/mRETjzFCn8eQ4wTaVn0DVI5fDrzHQkWJZGwXGT1jHd3kgIhR
vnnt4/s1GS4y90iqr9h3uXogUiFnrvHkgefZFMyUR3b9g2C58V5bCxrzKnIA/Ir7loTmotSl3WLc
q2PCTRuVepdRdzAytR2tSZDbeN8T+e6LnvTwZqAc0J7iljG7IWe3G11QXZ6Q1xpqvoXhhCOa/vNc
8zAghC4xlT6uww826zV+aksXRcKKRmQpmTnagXZyZKfoi4AdrvxCPwUIvjfWwkB16OUzh4aK15eT
4hLuCXGZ6mYlDtFvZGGePSCP6ue5D5b7gDWlPECYULivqMtrnCCeqlq9yMNT3ZFHV5FNZnHqTrs0
jF0ps56H3rQ/VmnMXOTWz6jSlECa2FD4xTV/qva2tj/as6WEKwqjGjr5vXq4dop0OpS/PGZZHGvn
vaiPUDGzA2Fd3/V20HBf+vjRMJzaZAeY+IiFcC3+NEJ6PmvFODTCCxf+nyN7IYPE8n2oPkxG7GZu
NksZM5ZHKvggMa41EwOQXEflA0VbxVDznbBtrD7vbPRF44SU1tN0oOVvMnSgXv8eDiVTgnQPYCrR
obzVDOS8MffUYNtUOwvEm7nCjypXc8DjMP62fU2jc5ZwrClJvGNSxjRMFbVPY4qcbBii2YQfmWs9
QqRJErH/LWYw3MFWaRPhCaYhhNsb0sUn0/36eVnSqUnQTu1r9m+37OZhHzHWcISBRS4coT8RFwtg
96cusBAO6RycUwPQWoa01kM2mbSgrhX9Z5+/Kh4604UO3ZqnleWphS22BtzMEopSvIdxrqID0Oqc
RnhLvbV/8a3hKpVO+n8+XbwYaLiuC3KZOixDvR0f4Fb4GiNAfpuRHAYr71rSFG1PPK0JsOivX3ZM
HtzQqKM//1s1apiKr1Bf/7xVCCb+5LHn70cUn3W9Onp5F0zCkZIACUcZQrbtG7obDm51m8YV/FoR
MpXLiBqAh5uhvcTGNQ6KZ4qQhJBGQAsRKl/TSXUHcDsYfJimh/u/VLjXmygK5M/cYw2k2gIp0GD2
q+a0CSg5lJMTuqgEeDC+wFgvQsfILOSB2NpE6EOXxvQrfFWUzktAIbSiKVJ9wPcboYqWevbCIiKt
irQfS2cfXeKi81bTzhQH5x3Y1ikx4+5ncBQUfXBoMVOmee8ipTLZcfxb0dp7BGOwj3pdBBc4jPWs
+Ecg6f5Eg9wegqMfaXqBLtME56S6c3/u/rk36s0WEuPfSgdf4sT/LKkH6XekJZJ0wCyz9FPTK1J2
D+NBda93rfmMOvplyEez10Zzh6bO1+jwC2joE3qAfKnCBnlKCFuM+NIMwdMSS2QZu1kxKMrejML5
3rqcp6iKIb8iAdvK/tCxbO6srOda7WFPg+TB/y2Wab5BWdTh0VFm3AI1Hv75jwfoePE2t4QOu9nH
d+1E/7bk3QA4DU6w1oxREfW5KdBHf78/XDKfTAJqWxAYF4irpwWsnWHvGpptsul8gyfD2koWPSSH
QRNy8nPMr1Kk9tE38eCXg5osk4XaGvArlvNbQL+f44S1F/r07WSiTGN0xgXF/WM0WDePjN9DJb6/
2dzrqJR2xqsXII8P7xnSDqyef0RinFM68aGh6jblwJ9/S4v2ygBcnZqjP/pXU1bRX2T5X7+UaYtA
rZhtuekYGDMJ6Q7Dm82joJnmg4U9gFrzScH3DAOqJT28DK2aMHirtjGKebxLXOd+CKMunh8NZdZR
zfLqE4W7Tfd+nAdX9Sg9B99MYGby97ivl2AzHRu3P0/kAoScOvwCD074BMVTBOH/vF4wtix5Mbgh
SMtSzAcBX/Ksticc7/3F63rKxJDBHgCt+ChdtZNkGwYu4ksfWo8E39i3813d5fj61P/rEI1QzIF4
gKNkMg4oKsP1uQAE3SsrfQY8XVN0o/MAkWkbGixa2FmQNK03uga3GMgV5bPBC5q66XFAkGIVD7Nf
aVkrF1tvEXHIrX/MrIxOT83gtV6COFxkTgAxjLNHqf+NL91aB2H6NvDPx3DyrboRtonMAxEVdVN6
kDBqx4MDnoypUiP9wwKSZBKlXZ52fS74gJo7WBKiFdR8YXYqeAPGD+LYwliDhp7ek4vJlsT9IM1i
A9r1ForEi2YcOB3EiSvBYYniw8w3DUQKLVAdu85yLlgbtBuVaKZu0O886sbUC3HhlNuBmzgP5/v/
Hd8Irzzx+Qe2s8NgqWbq8I66Mfli2vD04GlYPjvBNr92PmZe3qzYwQZXP5mn4voECGCDrRVYZira
X9RAuEp3EDG38ommVxuatceghd90JXWEwze/BnPAeNY5a6gPIFRO2DPSLptKivWuJ0lfzSsXo6ek
+0EAKEasUa5Qcx3Q+4fwzm64PE96ek90slWNby6LDt3fJSbOOwWryWAWkjpx5DiuDbn5HA3NJC27
OPg/n37PD7dKhhRw5iaJQyAm2sxbuKnuBvXK8/4M2acAq65HTzppRg0EOA1TAX77UE/5LKVKK840
WKOEdguvqtyd02QV1K990jvvLmNyIqQgtkLHewzy6jTV7z5/Uquw0iUY9w4nDiOQGkYClwyf5DID
B/TEzfb5hZxTv+Mx8AMIqZXfCB6JUBAUHrh4uZHduKvSjoKppgQ9XWv9uXEFNndk2WLVle4CDpex
aJLOoGrF+PseSfwdoZDKoTij+Ep5WcAT3uN6DpW4ZzaJYkQmpKroVYnP9uINkttlPfbFq+UKrkXv
DLe7iQPPsZkeQd+y9jGEqPtx4cPh9LjJA1T5/MQ6vK4eJf6ZKxsXs9bS4rcDcYNRDNh7NFmt4eJH
IMMdlZ4OzFl4kGCxfk5Cdg055coym05WTFX42PPFlXoFHWz1D03k2PoX2zgc1sMjuIE0pVGJg5Mu
lnER5786bRHLRXz3xGCfLJnaGx5oMtX1MK3GkWAwsFElu4wiwBtjmihgHnPxJAGJb2y/2K1j+DQY
8TCFx87+LOCKcm99s5zQ4LgZvZ8MbvirsdXWyy3ei/tnvJKG4o0WyAEDuJJLyUGzqbEOhfkCi2Ac
vgdYu0LAHgHyTzLPKKrYLvnY+F7RPjdGFczmu9Q1hgS/0ou2WArsVuMdadzmCUoMdzvZKZrjkluJ
SltGLQKOGFps1ae0j3NpSuVrhsGgQTuT6kRq4gytCJ2X734t0jRC+4+MztWrVH9KKWn0qdNw7BOk
RNKNdwdYieZB7zJGQ9MidG4gz10MIg0HCJPmmeDNjPz9tUHx4vSHuz++ghigHVmngM2gaz2INgdd
XZBZZvG18mGyMJY0MT8xxBtC31tFKVXJ2R4ED8wVUcQo5fOn12c3Eloy4krTljkgHRgs5SvK/n7u
cT2fXOTfWwkVSgFmvqdLF4BHwns0gHGwjpgjouUeoNgfslvmwJjkvMo7vdA1AHXGovO0OCK+4eQM
j4F1qXWHNpW0rEUC6PU4PELnssOQQrNZHK9w6TWlKT7B1l90b0d2YKodW+R34NdZzJpsPL98Dr0g
mdfiotiRKRY1dEcddcddmf6nuQKrecuLMj+8LrRerflDCqm1cpvJByFZrTZcczjOsM+vMawvhCeW
fW8xtrH0HDi5wY7DNAWLcNrcUJZ+cEcOlR10JF/J2Fetfq0anNilgnwD2rAdXej41sPYD5y6PPHf
pXoPlH4clauJ1CQBsZqtQO6+rXV04VkYasamfDWxgxTQJQcwYXBt/WH01yO9Wx297Cq470cRT74R
N8UT3N7aW5/rO4IuwsKSV49jXoYt0VYHeG+O221bpcmgRwM+SRTnY5wIlJBBanEtkmctkTJIU9wL
C2Pd9KBb45rH35hFdX8ffdCrdtKkQ8Zfe9+nd+j3+SYSCex8MyXc3GLZVkQn7FVXlssS/B2g3tp8
efQAO2ywLXKL5SzwOTtGABcrSV4AT6zLBCCvFN5wkUQnkHA20ecEPvgY+V23gIMQFhKtZq9eezcD
bigxnPKboEoEfBezND4vnvKBNOQFnrpOMXTX2zkJPP4sybG2XvvagjO3FxTTRZxJJpalkiACKk/i
SnxEk2nERoNlGtxsbpHItKlpuWxcNMcpDZZsHk2ITJOWeC3d6Lxo/n0h6h4/xKJGL/c1p5qV2mja
doGxfTvIQ/pQex3BX7/YF6iSVbtP2PUcxgeWXzkjqKb8ENSFZjAyosLaSi9jhD19umDn9oOnmDe3
2EOIko0XluXF3tvSgbo6dsCviSSopl7Kg0AsWmbD/fopSuSBdBAUDqV0N/lPSdaYTQCZ4eXKbIGs
uoTeJ0ebgRdCl8tyW+PG4T/feynb+I5dtN+YT0exXC933duLL14FfGhgTOvcHRlz1PHkMasqvupA
0hBQTHhoC3P/+2z5gz4OHvWKxOIFLv8eiOAb8qK6ZpNcIe5wZZr1Fngddr7D+WqQJJ2hayDvuc0P
0WbjT0S5RQDbV2LANrhK+ygGNrP64HLxGlFC492L80rPN+WKBFw0RMbsd+ioN2cD+Omkz7D1LyVT
BH7qQEmf6WrnQokR8IHjeNsRtrgdU5UnfvfYZScMJhYJFYhqpDVwZOchg0+Y9NYY9uMHlfh1GicH
6FdSSBtiAULuldZwc/BC9ZMobJ8Kxg==
`protect end_protected
